//==============================================================================
// ldpcenc_tbl.v
//
// Tables for 12 cyclic shifters.
//------------------------------------------------------------------------------
// Copyright (c) 2019 Guangxi Liu
//
// This source code is licensed under the MIT license found in the
// LICENSE file in the root directory of this source tree.
//==============================================================================


module ldpcenc_tbl (
    // System signals
    input clk,                  // system clock

    // Data interface
    input [8:0] addr,           // read address, [4:0]:cnt, [6:5]:rate, [8:7]:codeword length
    output reg [7:0] sh1,       // shift number for RCS1
    output reg [7:0] sh2,       // shift number for RCS2
    output reg [7:0] sh3,       // shift number for RCS3
    output reg [7:0] sh4,       // shift number for RCS4
    output reg [7:0] sh5,       // shift number for RCS5
    output reg [7:0] sh6,       // shift number for RCS6
    output reg [7:0] sh7,       // shift number for RCS7
    output reg [7:0] sh8,       // shift number for RCS8
    output reg [7:0] sh9,       // shift number for RCS9
    output reg [7:0] sh10,      // shift number for RCS10
    output reg [7:0] sh11,      // shift number for RCS11
    output reg [7:0] sh12       // shift number for RCS12
);

// Local signals
reg [7:0] sh1_w;
reg [7:0] sh2_w;
reg [7:0] sh3_w;
reg [7:0] sh4_w;
reg [7:0] sh5_w;
reg [7:0] sh6_w;
reg [7:0] sh7_w;
reg [7:0] sh8_w;
reg [7:0] sh9_w;
reg [7:0] sh10_w;
reg [7:0] sh11_w;
reg [7:0] sh12_w;


// Tables
always @ (*) begin
    case (addr)
        9'b00_00_00000: sh1_w = 8'd128;
        9'b00_00_00100: sh1_w = 8'd128;
        9'b00_00_00101: sh1_w = 8'd128;
        9'b00_00_01000: sh1_w = 8'd128;
        9'b00_00_01011: sh1_w = 8'd128;
        9'b00_01_00000: sh1_w = 8'd153;
        9'b00_01_00001: sh1_w = 8'd154;
        9'b00_01_00010: sh1_w = 8'd142;
        9'b00_01_00100: sh1_w = 8'd148;
        9'b00_01_00110: sh1_w = 8'd130;
        9'b00_01_01000: sh1_w = 8'd132;
        9'b00_01_01011: sh1_w = 8'd136;
        9'b00_01_01101: sh1_w = 8'd144;
        9'b00_01_01111: sh1_w = 8'd146;
        9'b00_10_00000: sh1_w = 8'd144;
        9'b00_10_00001: sh1_w = 8'd145;
        9'b00_10_00010: sh1_w = 8'd150;
        9'b00_10_00011: sh1_w = 8'd152;
        9'b00_10_00100: sh1_w = 8'd137;
        9'b00_10_00101: sh1_w = 8'd131;
        9'b00_10_00110: sh1_w = 8'd142;
        9'b00_10_01000: sh1_w = 8'd132;
        9'b00_10_01001: sh1_w = 8'd130;
        9'b00_10_01010: sh1_w = 8'd135;
        9'b00_10_01100: sh1_w = 8'd154;
        9'b00_10_01110: sh1_w = 8'd130;
        9'b00_10_10000: sh1_w = 8'd149;
        9'b00_11_00000: sh1_w = 8'd145;
        9'b00_11_00001: sh1_w = 8'd141;
        9'b00_11_00010: sh1_w = 8'd136;
        9'b00_11_00011: sh1_w = 8'd149;
        9'b00_11_00100: sh1_w = 8'd137;
        9'b00_11_00101: sh1_w = 8'd131;
        9'b00_11_00110: sh1_w = 8'd146;
        9'b00_11_00111: sh1_w = 8'd140;
        9'b00_11_01000: sh1_w = 8'd138;
        9'b00_11_01001: sh1_w = 8'd128;
        9'b00_11_01010: sh1_w = 8'd132;
        9'b00_11_01011: sh1_w = 8'd143;
        9'b00_11_01100: sh1_w = 8'd147;
        9'b00_11_01101: sh1_w = 8'd130;
        9'b00_11_01110: sh1_w = 8'd133;
        9'b00_11_01111: sh1_w = 8'd138;
        9'b00_11_10000: sh1_w = 8'd154;
        9'b00_11_10001: sh1_w = 8'd147;
        9'b00_11_10010: sh1_w = 8'd141;
        9'b00_11_10011: sh1_w = 8'd141;
        9'b01_00_00000: sh1_w = 8'd168;
        9'b01_00_00100: sh1_w = 8'd150;
        9'b01_00_00110: sh1_w = 8'd177;
        9'b01_00_00111: sh1_w = 8'd151;
        9'b01_00_01000: sh1_w = 8'd171;
        9'b01_01_00000: sh1_w = 8'd167;
        9'b01_01_00001: sh1_w = 8'd159;
        9'b01_01_00010: sh1_w = 8'd150;
        9'b01_01_00011: sh1_w = 8'd171;
        9'b01_01_00101: sh1_w = 8'd168;
        9'b01_01_00110: sh1_w = 8'd132;
        9'b01_01_01000: sh1_w = 8'd139;
        9'b01_01_01011: sh1_w = 8'd178;
        9'b01_01_01111: sh1_w = 8'd134;
        9'b01_10_00000: sh1_w = 8'd167;
        9'b01_10_00001: sh1_w = 8'd168;
        9'b01_10_00010: sh1_w = 8'd179;
        9'b01_10_00011: sh1_w = 8'd169;
        9'b01_10_00100: sh1_w = 8'd131;
        9'b01_10_00101: sh1_w = 8'd157;
        9'b01_10_00110: sh1_w = 8'd136;
        9'b01_10_00111: sh1_w = 8'd164;
        9'b01_10_01001: sh1_w = 8'd142;
        9'b01_10_01011: sh1_w = 8'd134;
        9'b01_10_01101: sh1_w = 8'd161;
        9'b01_10_01111: sh1_w = 8'd139;
        9'b01_10_10001: sh1_w = 8'd132;
        9'b01_11_00000: sh1_w = 8'd176;
        9'b01_11_00001: sh1_w = 8'd157;
        9'b01_11_00010: sh1_w = 8'd165;
        9'b01_11_00011: sh1_w = 8'd180;
        9'b01_11_00100: sh1_w = 8'd130;
        9'b01_11_00101: sh1_w = 8'd144;
        9'b01_11_00110: sh1_w = 8'd134;
        9'b01_11_00111: sh1_w = 8'd142;
        9'b01_11_01000: sh1_w = 8'd181;
        9'b01_11_01001: sh1_w = 8'd159;
        9'b01_11_01010: sh1_w = 8'd162;
        9'b01_11_01011: sh1_w = 8'd133;
        9'b01_11_01100: sh1_w = 8'd146;
        9'b01_11_01101: sh1_w = 8'd170;
        9'b01_11_01110: sh1_w = 8'd181;
        9'b01_11_01111: sh1_w = 8'd159;
        9'b01_11_10000: sh1_w = 8'd173;
        9'b01_11_10010: sh1_w = 8'd174;
        9'b01_11_10011: sh1_w = 8'd180;
        9'b10_00_00000: sh1_w = 8'd185;
        9'b10_00_00100: sh1_w = 8'd178;
        9'b10_00_00110: sh1_w = 8'd139;
        9'b10_00_01000: sh1_w = 8'd178;
        9'b10_00_01010: sh1_w = 8'd207;
        9'b10_01_00000: sh1_w = 8'd189;
        9'b10_01_00001: sh1_w = 8'd203;
        9'b10_01_00010: sh1_w = 8'd132;
        9'b10_01_00011: sh1_w = 8'd191;
        9'b10_01_00100: sh1_w = 8'd184;
        9'b10_01_01011: sh1_w = 8'd136;
        9'b10_01_01101: sh1_w = 8'd130;
        9'b10_01_01110: sh1_w = 8'd145;
        9'b10_01_01111: sh1_w = 8'd153;
        9'b10_10_00000: sh1_w = 8'd176;
        9'b10_10_00001: sh1_w = 8'd157;
        9'b10_10_00010: sh1_w = 8'd156;
        9'b10_10_00011: sh1_w = 8'd167;
        9'b10_10_00100: sh1_w = 8'd137;
        9'b10_10_00101: sh1_w = 8'd189;
        9'b10_10_01001: sh1_w = 8'd191;
        9'b10_10_01010: sh1_w = 8'd173;
        9'b10_10_01011: sh1_w = 8'd208;
        9'b10_10_01111: sh1_w = 8'd165;
        9'b10_10_10000: sh1_w = 8'd160;
        9'b10_10_10001: sh1_w = 8'd150;
        9'b10_11_00000: sh1_w = 8'd141;
        9'b10_11_00001: sh1_w = 8'd176;
        9'b10_11_00010: sh1_w = 8'd208;
        9'b10_11_00011: sh1_w = 8'd194;
        9'b10_11_00100: sh1_w = 8'd132;
        9'b10_11_00101: sh1_w = 8'd202;
        9'b10_11_00110: sh1_w = 8'd135;
        9'b10_11_00111: sh1_w = 8'd158;
        9'b10_11_01000: sh1_w = 8'd204;
        9'b10_11_01001: sh1_w = 8'd180;
        9'b10_11_01010: sh1_w = 8'd165;
        9'b10_11_01011: sh1_w = 8'd188;
        9'b10_11_01101: sh1_w = 8'd177;
        9'b10_11_01110: sh1_w = 8'd201;
        9'b10_11_01111: sh1_w = 8'd159;
        9'b10_11_10000: sh1_w = 8'd202;
        9'b10_11_10001: sh1_w = 8'd201;
        9'b10_11_10010: sh1_w = 8'd151;
        default: sh1_w = 8'd0;
    endcase
end

always @ (*) begin
    case (addr)
        9'b00_00_00000: sh2_w = 8'd150;
        9'b00_00_00001: sh2_w = 8'd128;
        9'b00_00_00100: sh2_w = 8'd145;
        9'b00_00_00110: sh2_w = 8'd128;
        9'b00_00_00111: sh2_w = 8'd128;
        9'b00_00_01000: sh2_w = 8'd140;
        9'b00_01_00000: sh2_w = 8'd138;
        9'b00_01_00001: sh2_w = 8'd137;
        9'b00_01_00010: sh2_w = 8'd143;
        9'b00_01_00011: sh2_w = 8'd139;
        9'b00_01_00101: sh2_w = 8'd128;
        9'b00_01_00111: sh2_w = 8'd129;
        9'b00_01_01010: sh2_w = 8'd146;
        9'b00_01_01100: sh2_w = 8'd136;
        9'b00_01_01110: sh2_w = 8'd138;
        9'b00_10_00000: sh2_w = 8'd153;
        9'b00_10_00001: sh2_w = 8'd140;
        9'b00_10_00010: sh2_w = 8'd140;
        9'b00_10_00011: sh2_w = 8'd131;
        9'b00_10_00100: sh2_w = 8'd131;
        9'b00_10_00101: sh2_w = 8'd154;
        9'b00_10_00110: sh2_w = 8'd134;
        9'b00_10_00111: sh2_w = 8'd149;
        9'b00_10_01001: sh2_w = 8'd143;
        9'b00_10_01010: sh2_w = 8'd150;
        9'b00_10_01100: sh2_w = 8'd143;
        9'b00_10_01110: sh2_w = 8'd132;
        9'b00_10_10001: sh2_w = 8'd144;
        9'b00_11_00000: sh2_w = 8'd131;
        9'b00_11_00001: sh2_w = 8'd140;
        9'b00_11_00010: sh2_w = 8'd139;
        9'b00_11_00011: sh2_w = 8'd142;
        9'b00_11_00100: sh2_w = 8'd139;
        9'b00_11_00101: sh2_w = 8'd153;
        9'b00_11_00110: sh2_w = 8'd133;
        9'b00_11_00111: sh2_w = 8'd146;
        9'b00_11_01000: sh2_w = 8'd128;
        9'b00_11_01001: sh2_w = 8'd137;
        9'b00_11_01010: sh2_w = 8'd130;
        9'b00_11_01011: sh2_w = 8'd154;
        9'b00_11_01100: sh2_w = 8'd154;
        9'b00_11_01101: sh2_w = 8'd138;
        9'b00_11_01110: sh2_w = 8'd152;
        9'b00_11_01111: sh2_w = 8'd135;
        9'b00_11_10000: sh2_w = 8'd142;
        9'b00_11_10001: sh2_w = 8'd148;
        9'b00_11_10010: sh2_w = 8'd132;
        9'b00_11_10011: sh2_w = 8'd130;
        9'b01_00_00000: sh2_w = 8'd178;
        9'b01_00_00001: sh2_w = 8'd129;
        9'b01_00_00100: sh2_w = 8'd176;
        9'b01_00_00101: sh2_w = 8'd163;
        9'b01_00_01000: sh2_w = 8'd141;
        9'b01_00_01010: sh2_w = 8'd158;
        9'b01_01_00000: sh2_w = 8'd153;
        9'b01_01_00001: sh2_w = 8'd180;
        9'b01_01_00010: sh2_w = 8'd169;
        9'b01_01_00011: sh2_w = 8'd130;
        9'b01_01_00100: sh2_w = 8'd134;
        9'b01_01_00110: sh2_w = 8'd142;
        9'b01_01_01000: sh2_w = 8'd162;
        9'b01_01_01100: sh2_w = 8'd152;
        9'b01_01_01110: sh2_w = 8'd165;
        9'b01_10_00000: sh2_w = 8'd176;
        9'b01_10_00001: sh2_w = 8'd149;
        9'b01_10_00010: sh2_w = 8'd175;
        9'b01_10_00011: sh2_w = 8'd137;
        9'b01_10_00100: sh2_w = 8'd176;
        9'b01_10_00101: sh2_w = 8'd163;
        9'b01_10_00110: sh2_w = 8'd179;
        9'b01_10_01000: sh2_w = 8'd166;
        9'b01_10_01010: sh2_w = 8'd156;
        9'b01_10_01100: sh2_w = 8'd162;
        9'b01_10_01110: sh2_w = 8'd178;
        9'b01_10_10000: sh2_w = 8'd178;
        9'b01_11_00000: sh2_w = 8'd145;
        9'b01_11_00001: sh2_w = 8'd132;
        9'b01_11_00010: sh2_w = 8'd158;
        9'b01_11_00011: sh2_w = 8'd135;
        9'b01_11_00100: sh2_w = 8'd171;
        9'b01_11_00101: sh2_w = 8'd139;
        9'b01_11_00110: sh2_w = 8'd152;
        9'b01_11_00111: sh2_w = 8'd134;
        9'b01_11_01000: sh2_w = 8'd142;
        9'b01_11_01001: sh2_w = 8'd149;
        9'b01_11_01010: sh2_w = 8'd134;
        9'b01_11_01011: sh2_w = 8'd167;
        9'b01_11_01100: sh2_w = 8'd145;
        9'b01_11_01101: sh2_w = 8'd168;
        9'b01_11_01110: sh2_w = 8'd175;
        9'b01_11_01111: sh2_w = 8'd135;
        9'b01_11_10000: sh2_w = 8'd143;
        9'b01_11_10001: sh2_w = 8'd169;
        9'b01_11_10010: sh2_w = 8'd147;
        9'b10_00_00000: sh2_w = 8'd131;
        9'b10_00_00010: sh2_w = 8'd156;
        9'b10_00_00100: sh2_w = 8'd128;
        9'b10_00_01000: sh2_w = 8'd183;
        9'b10_00_01001: sh2_w = 8'd135;
        9'b10_01_00000: sh2_w = 8'd184;
        9'b10_01_00001: sh2_w = 8'd202;
        9'b10_01_00010: sh2_w = 8'd205;
        9'b10_01_00011: sh2_w = 8'd148;
        9'b10_01_00111: sh2_w = 8'd192;
        9'b10_01_01000: sh2_w = 8'd152;
        9'b10_01_01001: sh2_w = 8'd132;
        9'b10_01_01010: sh2_w = 8'd195;
        9'b10_01_01100: sh2_w = 8'd135;
        9'b10_10_00000: sh2_w = 8'd132;
        9'b10_10_00001: sh2_w = 8'd177;
        9'b10_10_00010: sh2_w = 8'd170;
        9'b10_10_00011: sh2_w = 8'd176;
        9'b10_10_00100: sh2_w = 8'd139;
        9'b10_10_00101: sh2_w = 8'd158;
        9'b10_10_01001: sh2_w = 8'd177;
        9'b10_10_01010: sh2_w = 8'd145;
        9'b10_10_01011: sh2_w = 8'd169;
        9'b10_10_01100: sh2_w = 8'd165;
        9'b10_10_01101: sh2_w = 8'd143;
        9'b10_10_01111: sh2_w = 8'd182;
        9'b10_11_00000: sh2_w = 8'd197;
        9'b10_11_00001: sh2_w = 8'd191;
        9'b10_11_00010: sh2_w = 8'd202;
        9'b10_11_00011: sh2_w = 8'd184;
        9'b10_11_00100: sh2_w = 8'd192;
        9'b10_11_00101: sh2_w = 8'd205;
        9'b10_11_00110: sh2_w = 8'd185;
        9'b10_11_00111: sh2_w = 8'd193;
        9'b10_11_01000: sh2_w = 8'd134;
        9'b10_11_01001: sh2_w = 8'd144;
        9'b10_11_01010: sh2_w = 8'd179;
        9'b10_11_01100: sh2_w = 8'd192;
        9'b10_11_01110: sh2_w = 8'd196;
        9'b10_11_01111: sh2_w = 8'd137;
        9'b10_11_10000: sh2_w = 8'd176;
        9'b10_11_10001: sh2_w = 8'd190;
        9'b10_11_10010: sh2_w = 8'd182;
        9'b10_11_10011: sh2_w = 8'd155;
        default: sh2_w = 8'd0;
    endcase
end

always @ (*) begin
    case (addr)
        9'b00_00_00000: sh3_w = 8'd134;
        9'b00_00_00010: sh3_w = 8'd128;
        9'b00_00_00100: sh3_w = 8'd138;
        9'b00_00_01000: sh3_w = 8'd152;
        9'b00_00_01010: sh3_w = 8'd128;
        9'b00_01_00000: sh3_w = 8'd144;
        9'b00_01_00001: sh3_w = 8'd130;
        9'b00_01_00010: sh3_w = 8'd148;
        9'b00_01_00011: sh3_w = 8'd154;
        9'b00_01_00100: sh3_w = 8'd149;
        9'b00_01_00110: sh3_w = 8'd134;
        9'b00_01_01000: sh3_w = 8'd129;
        9'b00_01_01001: sh3_w = 8'd154;
        9'b00_01_01011: sh3_w = 8'd135;
        9'b00_10_00000: sh3_w = 8'd153;
        9'b00_10_00001: sh3_w = 8'd146;
        9'b00_10_00010: sh3_w = 8'd154;
        9'b00_10_00011: sh3_w = 8'd144;
        9'b00_10_00100: sh3_w = 8'd150;
        9'b00_10_00101: sh3_w = 8'd151;
        9'b00_10_00110: sh3_w = 8'd137;
        9'b00_10_01000: sh3_w = 8'd128;
        9'b00_10_01010: sh3_w = 8'd132;
        9'b00_10_01100: sh3_w = 8'd132;
        9'b00_10_01110: sh3_w = 8'd136;
        9'b00_10_01111: sh3_w = 8'd151;
        9'b00_10_10000: sh3_w = 8'd139;
        9'b00_11_00000: sh3_w = 8'd150;
        9'b00_11_00001: sh3_w = 8'd144;
        9'b00_11_00010: sh3_w = 8'd132;
        9'b00_11_00011: sh3_w = 8'd131;
        9'b00_11_00100: sh3_w = 8'd138;
        9'b00_11_00101: sh3_w = 8'd149;
        9'b00_11_00110: sh3_w = 8'd140;
        9'b00_11_00111: sh3_w = 8'd133;
        9'b00_11_01000: sh3_w = 8'd149;
        9'b00_11_01001: sh3_w = 8'd142;
        9'b00_11_01010: sh3_w = 8'd147;
        9'b00_11_01011: sh3_w = 8'd133;
        9'b00_11_01101: sh3_w = 8'd136;
        9'b00_11_01110: sh3_w = 8'd133;
        9'b00_11_01111: sh3_w = 8'd146;
        9'b00_11_10000: sh3_w = 8'd139;
        9'b00_11_10001: sh3_w = 8'd133;
        9'b00_11_10010: sh3_w = 8'd133;
        9'b00_11_10011: sh3_w = 8'd143;
        9'b01_00_00000: sh3_w = 8'd167;
        9'b01_00_00001: sh3_w = 8'd178;
        9'b01_00_00100: sh3_w = 8'd132;
        9'b01_00_00110: sh3_w = 8'd130;
        9'b01_00_01011: sh3_w = 8'd177;
        9'b01_01_00000: sh3_w = 8'd171;
        9'b01_01_00001: sh3_w = 8'd159;
        9'b01_01_00010: sh3_w = 8'd157;
        9'b01_01_00011: sh3_w = 8'd128;
        9'b01_01_00100: sh3_w = 8'd149;
        9'b01_01_00110: sh3_w = 8'd156;
        9'b01_01_01001: sh3_w = 8'd130;
        9'b01_01_01100: sh3_w = 8'd135;
        9'b01_01_01110: sh3_w = 8'd145;
        9'b01_10_00000: sh3_w = 8'd158;
        9'b01_10_00001: sh3_w = 8'd167;
        9'b01_10_00010: sh3_w = 8'd156;
        9'b01_10_00011: sh3_w = 8'd170;
        9'b01_10_00100: sh3_w = 8'd178;
        9'b01_10_00101: sh3_w = 8'd167;
        9'b01_10_00110: sh3_w = 8'd133;
        9'b01_10_00111: sh3_w = 8'd145;
        9'b01_10_01001: sh3_w = 8'd134;
        9'b01_10_01011: sh3_w = 8'd146;
        9'b01_10_01101: sh3_w = 8'd148;
        9'b01_10_01111: sh3_w = 8'd143;
        9'b01_10_10001: sh3_w = 8'd168;
        9'b01_11_00000: sh3_w = 8'd135;
        9'b01_11_00001: sh3_w = 8'd130;
        9'b01_11_00010: sh3_w = 8'd179;
        9'b01_11_00011: sh3_w = 8'd159;
        9'b01_11_00100: sh3_w = 8'd174;
        9'b01_11_00101: sh3_w = 8'd151;
        9'b01_11_00110: sh3_w = 8'd144;
        9'b01_11_00111: sh3_w = 8'd139;
        9'b01_11_01000: sh3_w = 8'd181;
        9'b01_11_01001: sh3_w = 8'd168;
        9'b01_11_01010: sh3_w = 8'd138;
        9'b01_11_01011: sh3_w = 8'd135;
        9'b01_11_01100: sh3_w = 8'd174;
        9'b01_11_01101: sh3_w = 8'd181;
        9'b01_11_01110: sh3_w = 8'd161;
        9'b01_11_01111: sh3_w = 8'd163;
        9'b01_11_10001: sh3_w = 8'd153;
        9'b01_11_10010: sh3_w = 8'd163;
        9'b01_11_10011: sh3_w = 8'd166;
        9'b10_00_00000: sh3_w = 8'd158;
        9'b10_00_00100: sh3_w = 8'd152;
        9'b10_00_00101: sh3_w = 8'd165;
        9'b10_00_01000: sh3_w = 8'd184;
        9'b10_00_01001: sh3_w = 8'd142;
        9'b10_01_00000: sh3_w = 8'd156;
        9'b10_01_00001: sh3_w = 8'd149;
        9'b10_01_00010: sh3_w = 8'd196;
        9'b10_01_00011: sh3_w = 8'd138;
        9'b10_01_00100: sh3_w = 8'd135;
        9'b10_01_00101: sh3_w = 8'd142;
        9'b10_01_00110: sh3_w = 8'd193;
        9'b10_01_01010: sh3_w = 8'd151;
        9'b10_01_01110: sh3_w = 8'd203;
        9'b10_10_00000: sh3_w = 8'd163;
        9'b10_10_00001: sh3_w = 8'd204;
        9'b10_10_00010: sh3_w = 8'd206;
        9'b10_10_00011: sh3_w = 8'd179;
        9'b10_10_00100: sh3_w = 8'd165;
        9'b10_10_00101: sh3_w = 8'd163;
        9'b10_10_00110: sh3_w = 8'd149;
        9'b10_10_01000: sh3_w = 8'd145;
        9'b10_10_01001: sh3_w = 8'd192;
        9'b10_10_01101: sh3_w = 8'd187;
        9'b10_10_01110: sh3_w = 8'd135;
        9'b10_10_10001: sh3_w = 8'd160;
        9'b10_11_00000: sh3_w = 8'd179;
        9'b10_11_00001: sh3_w = 8'd143;
        9'b10_11_00010: sh3_w = 8'd128;
        9'b10_11_00011: sh3_w = 8'd208;
        9'b10_11_00100: sh3_w = 8'd152;
        9'b10_11_00101: sh3_w = 8'd153;
        9'b10_11_00110: sh3_w = 8'd170;
        9'b10_11_00111: sh3_w = 8'd182;
        9'b10_11_01000: sh3_w = 8'd172;
        9'b10_11_01001: sh3_w = 8'd199;
        9'b10_11_01010: sh3_w = 8'd199;
        9'b10_11_01011: sh3_w = 8'd137;
        9'b10_11_01100: sh3_w = 8'd195;
        9'b10_11_01101: sh3_w = 8'd163;
        9'b10_11_01111: sh3_w = 8'd186;
        9'b10_11_10001: sh3_w = 8'd157;
        9'b10_11_10011: sh3_w = 8'd181;
        default: sh3_w = 8'd0;
    endcase
end

always @ (*) begin
    case (addr)
        9'b00_00_00000: sh4_w = 8'd130;
        9'b00_00_00011: sh4_w = 8'd128;
        9'b00_00_00100: sh4_w = 8'd148;
        9'b00_00_01000: sh4_w = 8'd153;
        9'b00_00_01001: sh4_w = 8'd128;
        9'b00_01_00000: sh4_w = 8'd138;
        9'b00_01_00001: sh4_w = 8'd141;
        9'b00_01_00010: sh4_w = 8'd133;
        9'b00_01_00011: sh4_w = 8'd128;
        9'b00_01_00101: sh4_w = 8'd131;
        9'b00_01_00111: sh4_w = 8'd135;
        9'b00_01_01010: sh4_w = 8'd154;
        9'b00_01_01101: sh4_w = 8'd141;
        9'b00_01_01111: sh4_w = 8'd144;
        9'b00_10_00000: sh4_w = 8'd137;
        9'b00_10_00001: sh4_w = 8'd135;
        9'b00_10_00010: sh4_w = 8'd128;
        9'b00_10_00011: sh4_w = 8'd129;
        9'b00_10_00100: sh4_w = 8'd145;
        9'b00_10_00111: sh4_w = 8'd135;
        9'b00_10_01000: sh4_w = 8'd131;
        9'b00_10_01010: sh4_w = 8'd131;
        9'b00_10_01011: sh4_w = 8'd151;
        9'b00_10_01101: sh4_w = 8'd144;
        9'b00_10_10000: sh4_w = 8'd149;
        9'b00_11_00000: sh4_w = 8'd135;
        9'b00_11_00001: sh4_w = 8'd135;
        9'b00_11_00010: sh4_w = 8'd142;
        9'b00_11_00011: sh4_w = 8'd142;
        9'b00_11_00100: sh4_w = 8'd132;
        9'b00_11_00101: sh4_w = 8'd144;
        9'b00_11_00110: sh4_w = 8'd144;
        9'b00_11_00111: sh4_w = 8'd152;
        9'b00_11_01000: sh4_w = 8'd152;
        9'b00_11_01001: sh4_w = 8'd138;
        9'b00_11_01010: sh4_w = 8'd129;
        9'b00_11_01011: sh4_w = 8'd135;
        9'b00_11_01100: sh4_w = 8'd143;
        9'b00_11_01101: sh4_w = 8'd134;
        9'b00_11_01110: sh4_w = 8'd138;
        9'b00_11_01111: sh4_w = 8'd154;
        9'b00_11_10000: sh4_w = 8'd136;
        9'b00_11_10001: sh4_w = 8'd146;
        9'b00_11_10010: sh4_w = 8'd149;
        9'b00_11_10011: sh4_w = 8'd142;
        9'b01_00_00000: sh4_w = 8'd161;
        9'b01_00_00011: sh4_w = 8'd166;
        9'b01_00_00100: sh4_w = 8'd165;
        9'b01_00_00111: sh4_w = 8'd132;
        9'b01_00_01000: sh4_w = 8'd129;
        9'b01_01_00000: sh4_w = 8'd148;
        9'b01_01_00001: sh4_w = 8'd161;
        9'b01_01_00010: sh4_w = 8'd176;
        9'b01_01_00100: sh4_w = 8'd132;
        9'b01_01_00101: sh4_w = 8'd141;
        9'b01_01_00111: sh4_w = 8'd154;
        9'b01_01_01010: sh4_w = 8'd150;
        9'b01_01_01101: sh4_w = 8'd174;
        9'b01_01_01110: sh4_w = 8'd170;
        9'b01_10_00000: sh4_w = 8'd157;
        9'b01_10_00001: sh4_w = 8'd128;
        9'b01_10_00010: sh4_w = 8'd129;
        9'b01_10_00011: sh4_w = 8'd171;
        9'b01_10_00100: sh4_w = 8'd164;
        9'b01_10_00101: sh4_w = 8'd158;
        9'b01_10_00110: sh4_w = 8'd175;
        9'b01_10_01000: sh4_w = 8'd177;
        9'b01_10_01010: sh4_w = 8'd175;
        9'b01_10_01100: sh4_w = 8'd131;
        9'b01_10_01110: sh4_w = 8'd163;
        9'b01_10_10000: sh4_w = 8'd162;
        9'b01_11_00000: sh4_w = 8'd147;
        9'b01_11_00001: sh4_w = 8'd176;
        9'b01_11_00010: sh4_w = 8'd169;
        9'b01_11_00011: sh4_w = 8'd129;
        9'b01_11_00100: sh4_w = 8'd138;
        9'b01_11_00101: sh4_w = 8'd135;
        9'b01_11_00110: sh4_w = 8'd164;
        9'b01_11_00111: sh4_w = 8'd175;
        9'b01_11_01000: sh4_w = 8'd133;
        9'b01_11_01001: sh4_w = 8'd157;
        9'b01_11_01010: sh4_w = 8'd180;
        9'b01_11_01011: sh4_w = 8'd180;
        9'b01_11_01100: sh4_w = 8'd159;
        9'b01_11_01101: sh4_w = 8'd138;
        9'b01_11_01110: sh4_w = 8'd154;
        9'b01_11_01111: sh4_w = 8'd134;
        9'b01_11_10000: sh4_w = 8'd131;
        9'b01_11_10001: sh4_w = 8'd130;
        9'b01_11_10011: sh4_w = 8'd179;
        9'b10_00_00000: sh4_w = 8'd190;
        9'b10_00_00001: sh4_w = 8'd181;
        9'b10_00_00100: sh4_w = 8'd181;
        9'b10_00_00111: sh4_w = 8'd131;
        9'b10_00_01000: sh4_w = 8'd163;
        9'b10_01_00000: sh4_w = 8'd176;
        9'b10_01_00001: sh4_w = 8'd166;
        9'b10_01_00010: sh4_w = 8'd171;
        9'b10_01_00011: sh4_w = 8'd206;
        9'b10_01_00100: sh4_w = 8'd204;
        9'b10_01_01001: sh4_w = 8'd133;
        9'b10_01_01010: sh4_w = 8'd164;
        9'b10_01_01100: sh4_w = 8'd143;
        9'b10_01_01101: sh4_w = 8'd200;
        9'b10_10_00000: sh4_w = 8'd137;
        9'b10_10_00001: sh4_w = 8'd193;
        9'b10_10_00010: sh4_w = 8'd172;
        9'b10_10_00011: sh4_w = 8'd137;
        9'b10_10_00100: sh4_w = 8'd182;
        9'b10_10_00101: sh4_w = 8'd184;
        9'b10_10_00110: sh4_w = 8'd201;
        9'b10_10_00111: sh4_w = 8'd162;
        9'b10_10_01000: sh4_w = 8'd170;
        9'b10_10_01100: sh4_w = 8'd163;
        9'b10_10_10000: sh4_w = 8'd174;
        9'b10_10_10001: sh4_w = 8'd167;
        9'b10_11_00000: sh4_w = 8'd144;
        9'b10_11_00001: sh4_w = 8'd157;
        9'b10_11_00010: sh4_w = 8'd164;
        9'b10_11_00011: sh4_w = 8'd169;
        9'b10_11_00100: sh4_w = 8'd172;
        9'b10_11_00101: sh4_w = 8'd184;
        9'b10_11_00110: sh4_w = 8'd187;
        9'b10_11_00111: sh4_w = 8'd165;
        9'b10_11_01000: sh4_w = 8'd178;
        9'b10_11_01001: sh4_w = 8'd152;
        9'b10_11_01011: sh4_w = 8'd193;
        9'b10_11_01100: sh4_w = 8'd132;
        9'b10_11_01101: sh4_w = 8'd193;
        9'b10_11_01110: sh4_w = 8'd180;
        9'b10_11_10000: sh4_w = 8'd132;
        9'b10_11_10010: sh4_w = 8'd201;
        9'b10_11_10011: sh4_w = 8'd180;
        default: sh4_w = 8'd0;
    endcase
end

always @ (*) begin
    case (addr)
        9'b00_00_00000: sh5_w = 8'd151;
        9'b00_00_00100: sh5_w = 8'd131;
        9'b00_00_01000: sh5_w = 8'd128;
        9'b00_00_01010: sh5_w = 8'd137;
        9'b00_00_01011: sh5_w = 8'd139;
        9'b00_01_00000: sh5_w = 8'd151;
        9'b00_01_00001: sh5_w = 8'd142;
        9'b00_01_00010: sh5_w = 8'd152;
        9'b00_01_00100: sh5_w = 8'd140;
        9'b00_01_00110: sh5_w = 8'd147;
        9'b00_01_01000: sh5_w = 8'd145;
        9'b00_01_01100: sh5_w = 8'd148;
        9'b00_01_01110: sh5_w = 8'd149;
        9'b00_10_00000: sh5_w = 8'd152;
        9'b00_10_00001: sh5_w = 8'd133;
        9'b00_10_00010: sh5_w = 8'd154;
        9'b00_10_00011: sh5_w = 8'd135;
        9'b00_10_00100: sh5_w = 8'd129;
        9'b00_10_00111: sh5_w = 8'd143;
        9'b00_10_01000: sh5_w = 8'd152;
        9'b00_10_01001: sh5_w = 8'd143;
        9'b00_10_01011: sh5_w = 8'd136;
        9'b00_10_01101: sh5_w = 8'd141;
        9'b00_10_01111: sh5_w = 8'd141;
        9'b00_10_10001: sh5_w = 8'd139;
        9'b01_00_00000: sh5_w = 8'd173;
        9'b01_00_00100: sh5_w = 8'd128;
        9'b01_00_00101: sh5_w = 8'd150;
        9'b01_00_01000: sh5_w = 8'd148;
        9'b01_00_01001: sh5_w = 8'd170;
        9'b01_01_00000: sh5_w = 8'd173;
        9'b01_01_00001: sh5_w = 8'd135;
        9'b01_01_00010: sh5_w = 8'd146;
        9'b01_01_00011: sh5_w = 8'd179;
        9'b01_01_00100: sh5_w = 8'd140;
        9'b01_01_00101: sh5_w = 8'd153;
        9'b01_01_01001: sh5_w = 8'd178;
        9'b01_01_01100: sh5_w = 8'd133;
        9'b01_10_00000: sh5_w = 8'd129;
        9'b01_10_00001: sh5_w = 8'd160;
        9'b01_10_00010: sh5_w = 8'd139;
        9'b01_10_00011: sh5_w = 8'd151;
        9'b01_10_00100: sh5_w = 8'd138;
        9'b01_10_00101: sh5_w = 8'd172;
        9'b01_10_00110: sh5_w = 8'd140;
        9'b01_10_00111: sh5_w = 8'd135;
        9'b01_10_01001: sh5_w = 8'd176;
        9'b01_10_01011: sh5_w = 8'd132;
        9'b01_10_01101: sh5_w = 8'd137;
        9'b01_10_01111: sh5_w = 8'd145;
        9'b01_10_10001: sh5_w = 8'd144;
        9'b10_00_00000: sh5_w = 8'd168;
        9'b10_00_00011: sh5_w = 8'd148;
        9'b10_00_00100: sh5_w = 8'd194;
        9'b10_00_00111: sh5_w = 8'd150;
        9'b10_00_01000: sh5_w = 8'd156;
        9'b10_01_00000: sh5_w = 8'd168;
        9'b10_01_00001: sh5_w = 8'd130;
        9'b10_01_00010: sh5_w = 8'd181;
        9'b10_01_00011: sh5_w = 8'd153;
        9'b10_01_00101: sh5_w = 8'd180;
        9'b10_01_00110: sh5_w = 8'd190;
        9'b10_01_01000: sh5_w = 8'd148;
        9'b10_01_01011: sh5_w = 8'd172;
        9'b10_10_00000: sh5_w = 8'd131;
        9'b10_10_00001: sh5_w = 8'd190;
        9'b10_10_00010: sh5_w = 8'd135;
        9'b10_10_00011: sh5_w = 8'd208;
        9'b10_10_00100: sh5_w = 8'd196;
        9'b10_10_00101: sh5_w = 8'd154;
        9'b10_10_00111: sh5_w = 8'd208;
        9'b10_10_01000: sh5_w = 8'd183;
        9'b10_10_01010: sh5_w = 8'd164;
        9'b10_10_01100: sh5_w = 8'd154;
        9'b10_10_01110: sh5_w = 8'd137;
        9'b10_10_10000: sh5_w = 8'd200;
        default: sh5_w = 8'd0;
    endcase
end

always @ (*) begin
    case (addr)
        9'b00_00_00000: sh6_w = 8'd152;
        9'b00_00_00010: sh6_w = 8'd151;
        9'b00_00_00011: sh6_w = 8'd129;
        9'b00_00_00100: sh6_w = 8'd145;
        9'b00_00_00110: sh6_w = 8'd131;
        9'b00_00_01000: sh6_w = 8'd138;
        9'b00_01_00000: sh6_w = 8'd134;
        9'b00_01_00001: sh6_w = 8'd150;
        9'b00_01_00010: sh6_w = 8'd137;
        9'b00_01_00011: sh6_w = 8'd148;
        9'b00_01_00101: sh6_w = 8'd153;
        9'b00_01_00111: sh6_w = 8'd145;
        9'b00_01_01001: sh6_w = 8'd136;
        9'b00_01_01011: sh6_w = 8'd142;
        9'b00_01_01101: sh6_w = 8'd146;
        9'b00_10_00000: sh6_w = 8'd130;
        9'b00_10_00001: sh6_w = 8'd130;
        9'b00_10_00010: sh6_w = 8'd147;
        9'b00_10_00011: sh6_w = 8'd142;
        9'b00_10_00100: sh6_w = 8'd152;
        9'b00_10_00101: sh6_w = 8'd129;
        9'b00_10_00110: sh6_w = 8'd143;
        9'b00_10_00111: sh6_w = 8'd147;
        9'b00_10_01001: sh6_w = 8'd149;
        9'b00_10_01011: sh6_w = 8'd130;
        9'b00_10_01101: sh6_w = 8'd152;
        9'b00_10_01111: sh6_w = 8'd131;
        9'b00_10_10001: sh6_w = 8'd130;
        9'b01_00_00000: sh6_w = 8'd179;
        9'b01_00_00011: sh6_w = 8'd176;
        9'b01_00_00100: sh6_w = 8'd163;
        9'b01_00_01000: sh6_w = 8'd172;
        9'b01_00_01010: sh6_w = 8'd146;
        9'b01_01_00000: sh6_w = 8'd163;
        9'b01_01_00001: sh6_w = 8'd168;
        9'b01_01_00010: sh6_w = 8'd160;
        9'b01_01_00011: sh6_w = 8'd144;
        9'b01_01_00100: sh6_w = 8'd133;
        9'b01_01_00111: sh6_w = 8'd146;
        9'b01_01_01010: sh6_w = 8'd171;
        9'b01_01_01011: sh6_w = 8'd179;
        9'b01_01_01101: sh6_w = 8'd160;
        9'b01_10_00000: sh6_w = 8'd141;
        9'b01_10_00001: sh6_w = 8'd135;
        9'b01_10_00010: sh6_w = 8'd143;
        9'b01_10_00011: sh6_w = 8'd175;
        9'b01_10_00100: sh6_w = 8'd151;
        9'b01_10_00101: sh6_w = 8'd144;
        9'b01_10_00110: sh6_w = 8'd175;
        9'b01_10_01000: sh6_w = 8'd171;
        9'b01_10_01010: sh6_w = 8'd157;
        9'b01_10_01100: sh6_w = 8'd180;
        9'b01_10_01110: sh6_w = 8'd130;
        9'b01_10_10000: sh6_w = 8'd181;
        9'b10_00_00000: sh6_w = 8'd128;
        9'b10_00_00100: sh6_w = 8'd136;
        9'b10_00_00110: sh6_w = 8'd170;
        9'b10_00_01000: sh6_w = 8'd178;
        9'b10_00_01011: sh6_w = 8'd136;
        9'b10_01_00000: sh6_w = 8'd197;
        9'b10_01_00001: sh6_w = 8'd151;
        9'b10_01_00010: sh6_w = 8'd192;
        9'b10_01_00011: sh6_w = 8'd138;
        9'b10_01_00100: sh6_w = 8'd150;
        9'b10_01_00110: sh6_w = 8'd149;
        9'b10_01_01100: sh6_w = 8'd196;
        9'b10_01_01101: sh6_w = 8'd151;
        9'b10_01_01110: sh6_w = 8'd157;
        9'b10_10_00000: sh6_w = 8'd154;
        9'b10_10_00001: sh6_w = 8'd203;
        9'b10_10_00010: sh6_w = 8'd161;
        9'b10_10_00011: sh6_w = 8'd149;
        9'b10_10_00100: sh6_w = 8'd197;
        9'b10_10_00101: sh6_w = 8'd187;
        9'b10_10_00110: sh6_w = 8'd131;
        9'b10_10_00111: sh6_w = 8'd166;
        9'b10_10_01011: sh6_w = 8'd163;
        9'b10_10_01101: sh6_w = 8'd190;
        9'b10_10_01110: sh6_w = 8'd164;
        9'b10_10_01111: sh6_w = 8'd154;
        default: sh6_w = 8'd0;
    endcase
end

always @ (*) begin
    case (addr)
        9'b00_00_00000: sh7_w = 8'd153;
        9'b00_00_00100: sh7_w = 8'd136;
        9'b00_00_01000: sh7_w = 8'd135;
        9'b00_00_01001: sh7_w = 8'd146;
        9'b00_01_00000: sh7_w = 8'd142;
        9'b00_01_00001: sh7_w = 8'd151;
        9'b00_01_00010: sh7_w = 8'd149;
        9'b00_01_00011: sh7_w = 8'd139;
        9'b00_01_00100: sh7_w = 8'd148;
        9'b00_01_00110: sh7_w = 8'd152;
        9'b00_01_01000: sh7_w = 8'd146;
        9'b00_01_01010: sh7_w = 8'd147;
        9'b00_01_01111: sh7_w = 8'd150;
        9'b01_00_00000: sh7_w = 8'd175;
        9'b01_00_00001: sh7_w = 8'd139;
        9'b01_00_00101: sh7_w = 8'd145;
        9'b01_00_01000: sh7_w = 8'd179;
        9'b01_01_00000: sh7_w = 8'd137;
        9'b01_01_00001: sh7_w = 8'd152;
        9'b01_01_00010: sh7_w = 8'd141;
        9'b01_01_00011: sh7_w = 8'd150;
        9'b01_01_00100: sh7_w = 8'd156;
        9'b01_01_00111: sh7_w = 8'd165;
        9'b01_01_01010: sh7_w = 8'd153;
        9'b01_01_01101: sh7_w = 8'd180;
        9'b01_01_01111: sh7_w = 8'd141;
        9'b10_00_00000: sh7_w = 8'd197;
        9'b10_00_00001: sh7_w = 8'd207;
        9'b10_00_00010: sh7_w = 8'd207;
        9'b10_00_00110: sh7_w = 8'd184;
        9'b10_00_01000: sh7_w = 8'd180;
        9'b10_01_00000: sh7_w = 8'd140;
        9'b10_01_00001: sh7_w = 8'd128;
        9'b10_01_00010: sh7_w = 8'd196;
        9'b10_01_00011: sh7_w = 8'd148;
        9'b10_01_00100: sh7_w = 8'd183;
        9'b10_01_00101: sh7_w = 8'd189;
        9'b10_01_00111: sh7_w = 8'd168;
        9'b10_01_01011: sh7_w = 8'd180;
        9'b10_01_01111: sh7_w = 8'd172;
        default: sh7_w = 8'd0;
    endcase
end

always @ (*) begin
    case (addr)
        9'b00_00_00000: sh8_w = 8'd141;
        9'b00_00_00001: sh8_w = 8'd152;
        9'b00_00_00100: sh8_w = 8'd128;
        9'b00_00_00110: sh8_w = 8'd136;
        9'b00_00_01000: sh8_w = 8'd134;
        9'b00_01_00000: sh8_w = 8'd145;
        9'b00_01_00001: sh8_w = 8'd139;
        9'b00_01_00010: sh8_w = 8'd139;
        9'b00_01_00011: sh8_w = 8'd148;
        9'b00_01_00101: sh8_w = 8'd149;
        9'b00_01_00111: sh8_w = 8'd154;
        9'b00_01_01001: sh8_w = 8'd131;
        9'b00_01_01100: sh8_w = 8'd146;
        9'b00_01_01110: sh8_w = 8'd154;
        9'b01_00_00000: sh8_w = 8'd133;
        9'b01_00_00010: sh8_w = 8'd153;
        9'b01_00_00100: sh8_w = 8'd134;
        9'b01_00_00110: sh8_w = 8'd173;
        9'b01_00_01000: sh8_w = 8'd141;
        9'b01_00_01001: sh8_w = 8'd168;
        9'b01_01_00000: sh8_w = 8'd160;
        9'b01_01_00001: sh8_w = 8'd150;
        9'b01_01_00010: sh8_w = 8'd132;
        9'b01_01_00011: sh8_w = 8'd149;
        9'b01_01_00100: sh8_w = 8'd144;
        9'b01_01_01000: sh8_w = 8'd155;
        9'b01_01_01001: sh8_w = 8'd156;
        9'b01_01_01011: sh8_w = 8'd166;
        9'b01_01_01111: sh8_w = 8'd136;
        9'b10_00_00000: sh8_w = 8'd193;
        9'b10_00_00100: sh8_w = 8'd166;
        9'b10_00_00101: sh8_w = 8'd185;
        9'b10_00_01000: sh8_w = 8'd200;
        9'b10_00_01010: sh8_w = 8'd155;
        9'b10_01_00000: sh8_w = 8'd186;
        9'b10_01_00001: sh8_w = 8'd136;
        9'b10_01_00010: sh8_w = 8'd162;
        9'b10_01_00011: sh8_w = 8'd192;
        9'b10_01_00100: sh8_w = 8'd206;
        9'b10_01_00111: sh8_w = 8'd139;
        9'b10_01_01000: sh8_w = 8'd206;
        9'b10_01_01001: sh8_w = 8'd152;
        9'b10_01_01111: sh8_w = 8'd186;
        default: sh8_w = 8'd0;
    endcase
end

always @ (*) begin
    case (addr)
        9'b00_00_00000: sh9_w = 8'd135;
        9'b00_00_00001: sh9_w = 8'd148;
        9'b00_00_00011: sh9_w = 8'd144;
        9'b00_00_00100: sh9_w = 8'd150;
        9'b00_00_00101: sh9_w = 8'd138;
        9'b00_00_01000: sh9_w = 8'd151;
        9'b01_00_00000: sh9_w = 8'd161;
        9'b01_00_00011: sh9_w = 8'd162;
        9'b01_00_00100: sh9_w = 8'd152;
        9'b01_00_01000: sh9_w = 8'd151;
        9'b01_00_01011: sh9_w = 8'd174;
        9'b10_00_00000: sh9_w = 8'd192;
        9'b10_00_00100: sh9_w = 8'd142;
        9'b10_00_00101: sh9_w = 8'd180;
        9'b10_00_01000: sh9_w = 8'd158;
        9'b10_00_01011: sh9_w = 8'd160;
        default: sh9_w = 8'd0;
    endcase
end

always @ (*) begin
    case (addr)
        9'b00_00_00000: sh10_w = 8'd139;
        9'b00_00_00100: sh10_w = 8'd147;
        9'b00_00_01000: sh10_w = 8'd141;
        9'b00_00_01010: sh10_w = 8'd131;
        9'b00_00_01011: sh10_w = 8'd145;
        9'b01_00_00000: sh10_w = 8'd129;
        9'b01_00_00010: sh10_w = 8'd155;
        9'b01_00_00100: sh10_w = 8'd129;
        9'b01_00_01000: sh10_w = 8'd166;
        9'b01_00_01010: sh10_w = 8'd172;
        9'b10_00_00001: sh10_w = 8'd173;
        9'b10_00_00011: sh10_w = 8'd198;
        9'b10_00_00100: sh10_w = 8'd128;
        9'b10_00_01000: sh10_w = 8'd205;
        9'b10_00_01001: sh10_w = 8'd137;
        default: sh10_w = 8'd0;
    endcase
end

always @ (*) begin
    case (addr)
        9'b00_00_00000: sh11_w = 8'd153;
        9'b00_00_00010: sh11_w = 8'd136;
        9'b00_00_00100: sh11_w = 8'd151;
        9'b00_00_00101: sh11_w = 8'd146;
        9'b00_00_00111: sh11_w = 8'd142;
        9'b00_00_01000: sh11_w = 8'd137;
        9'b01_00_00001: sh11_w = 8'd146;
        9'b01_00_00100: sh11_w = 8'd151;
        9'b01_00_00111: sh11_w = 8'd136;
        9'b01_00_01000: sh11_w = 8'd128;
        9'b01_00_01001: sh11_w = 8'd163;
        9'b10_00_00000: sh11_w = 8'd130;
        9'b10_00_00001: sh11_w = 8'd184;
        9'b10_00_00011: sh11_w = 8'd185;
        9'b10_00_00100: sh11_w = 8'd163;
        9'b10_00_01010: sh11_w = 8'd140;
        default: sh11_w = 8'd0;
    endcase
end

always @ (*) begin
    case (addr)
        9'b00_00_00000: sh12_w = 8'd131;
        9'b00_00_00100: sh12_w = 8'd144;
        9'b00_00_00111: sh12_w = 8'd130;
        9'b00_00_01000: sh12_w = 8'd153;
        9'b00_00_01001: sh12_w = 8'd133;
        9'b01_00_00000: sh12_w = 8'd177;
        9'b01_00_00010: sh12_w = 8'd145;
        9'b01_00_00100: sh12_w = 8'd158;
        9'b01_00_01000: sh12_w = 8'd162;
        9'b01_00_01011: sh12_w = 8'd147;
        9'b10_00_00000: sh12_w = 8'd152;
        9'b10_00_00010: sh12_w = 8'd189;
        9'b10_00_00100: sh12_w = 8'd188;
        9'b10_00_00111: sh12_w = 8'd155;
        9'b10_00_01000: sh12_w = 8'd179;
        9'b10_00_01011: sh12_w = 8'd144;
        default: sh12_w = 8'd0;
    endcase
end


// output data
always @ (posedge clk) begin
    sh1 <= sh1_w;
    sh2 <= sh2_w;
    sh3 <= sh3_w;
    sh4 <= sh4_w;
    sh5 <= sh5_w;
    sh6 <= sh6_w;
    sh7 <= sh7_w;
    sh8 <= sh8_w;
    sh9 <= sh9_w;
    sh10 <= sh10_w;
    sh11 <= sh11_w;
    sh12 <= sh12_w;
end


endmodule
